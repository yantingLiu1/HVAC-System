library ieee;
use ieee.std_logic_1164.all;

entity PB_Inverters is

	port(
		pb_in : IN std_logic_vector(3 downto 0);
		pb: out std_logic_vector(3 downto 0)
	);

end PB_Inverters;

architecture inverter of PB_Inverters is

	begin
	pb <= not(pb_in);

end inverter;